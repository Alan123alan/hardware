module Or(output out, input i1, input i0);
//modelling the circuit
or(out,i1,i0);
endmodule
