module mux_16_tb;
initial begin
$
end
endmodule
