module Not(input i0, output out);
//modeling the circuit
not(out, i0);
endmodule
