module And(output out, input i1, input i0);
// Modeling the circuit
and(out,i0,i1);
endmodule
