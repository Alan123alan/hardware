module SRLatch();
endmodule
