`include "../gates/Not16.v"
`include "../gates/And16.v"
`include "../demultiplexors/And16.v"
module ALU(output [15:0] out, input zx,nx,zy,ny,f,no, input [15:0] x, input [15:0] y);

endmodule
