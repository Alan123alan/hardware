module Mux4Way16(input [15:0] i0, input [15:0] i1, input [15:0] i2, input [15:0] i3, output [15:0] o);

endmodule
